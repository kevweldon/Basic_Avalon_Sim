// my_sys_reset_in.v

// Generated using ACDS version 23.4 79

`timescale 1 ps / 1 ps
module my_sys_reset_in (
		input  wire  clk,       //       clk.clk
		input  wire  in_reset,  //  in_reset.reset
		output wire  out_reset  // out_reset.reset
	);

	assign out_reset = in_reset;

endmodule
