// my_sys_clock_in.v

// Generated using ACDS version 23.1 115

`timescale 1 ps / 1 ps
module my_sys_clock_in (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);

	assign out_clk = in_clk;

endmodule
